VERSION 5.8 ;
BUSBITCHARS "[]" ;
DIVIDERCHAR "/" ;
UNITS
    DATABASE MICRONS 2000 ;
END UNITS
MACRO efuse_ctrl
  FOREIGN efuse_ctrl 0 0 ;
  CLASS BLOCK ;
  SIZE 2175 BY 2352.3 ;
  PIN wb_ack_o
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT  1887.2 0 1887.76 4 ;
    END
  END wb_ack_o
  PIN wb_adr_i[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT  39.2 0 39.76 4 ;
    END
  END wb_adr_i[0]
  PIN wb_adr_i[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT  655.2 0 655.76 4 ;
    END
  END wb_adr_i[10]
  PIN wb_adr_i[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT  716.8 0 717.36 4 ;
    END
  END wb_adr_i[11]
  PIN wb_adr_i[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT  100.8 0 101.36 4 ;
    END
  END wb_adr_i[1]
  PIN wb_adr_i[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT  162.4 0 162.96 4 ;
    END
  END wb_adr_i[2]
  PIN wb_adr_i[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT  224 0 224.56 4 ;
    END
  END wb_adr_i[3]
  PIN wb_adr_i[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT  285.6 0 286.16 4 ;
    END
  END wb_adr_i[4]
  PIN wb_adr_i[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT  347.2 0 347.76 4 ;
    END
  END wb_adr_i[5]
  PIN wb_adr_i[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT  408.8 0 409.36 4 ;
    END
  END wb_adr_i[6]
  PIN wb_adr_i[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT  470.4 0 470.96 4 ;
    END
  END wb_adr_i[7]
  PIN wb_adr_i[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT  532 0 532.56 4 ;
    END
  END wb_adr_i[8]
  PIN wb_adr_i[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT  593.6 0 594.16 4 ;
    END
  END wb_adr_i[9]
  PIN wb_clk_i
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT  2072 0 2072.56 4 ;
    END
  END wb_clk_i
  PIN wb_cyc_i
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT  2010.4 0 2010.96 4 ;
    END
  END wb_cyc_i
  PIN wb_dat_i[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT  1271.2 0 1271.76 4 ;
    END
  END wb_dat_i[0]
  PIN wb_dat_i[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT  1332.8 0 1333.36 4 ;
    END
  END wb_dat_i[1]
  PIN wb_dat_i[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT  1394.4 0 1394.96 4 ;
    END
  END wb_dat_i[2]
  PIN wb_dat_i[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT  1456 0 1456.56 4 ;
    END
  END wb_dat_i[3]
  PIN wb_dat_i[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT  1517.6 0 1518.16 4 ;
    END
  END wb_dat_i[4]
  PIN wb_dat_i[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT  1579.2 0 1579.76 4 ;
    END
  END wb_dat_i[5]
  PIN wb_dat_i[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT  1640.8 0 1641.36 4 ;
    END
  END wb_dat_i[6]
  PIN wb_dat_i[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT  1702.4 0 1702.96 4 ;
    END
  END wb_dat_i[7]
  PIN wb_dat_o[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT  778.4 0 778.96 4 ;
    END
  END wb_dat_o[0]
  PIN wb_dat_o[1]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT  840 0 840.56 4 ;
    END
  END wb_dat_o[1]
  PIN wb_dat_o[2]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT  901.6 0 902.16 4 ;
    END
  END wb_dat_o[2]
  PIN wb_dat_o[3]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT  963.2 0 963.76 4 ;
    END
  END wb_dat_o[3]
  PIN wb_dat_o[4]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT  1024.8 0 1025.36 4 ;
    END
  END wb_dat_o[4]
  PIN wb_dat_o[5]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT  1086.4 0 1086.96 4 ;
    END
  END wb_dat_o[5]
  PIN wb_dat_o[6]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT  1148 0 1148.56 4 ;
    END
  END wb_dat_o[6]
  PIN wb_dat_o[7]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT  1209.6 0 1210.16 4 ;
    END
  END wb_dat_o[7]
  PIN wb_rst_i
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT  2133.6 0 2134.16 4 ;
    END
  END wb_rst_i
  PIN wb_sel_i
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT  1948.8 0 1949.36 4 ;
    END
  END wb_sel_i
  PIN wb_stb_i
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT  1825.6 0 1826.16 4 ;
    END
  END wb_stb_i
  PIN wb_we_i
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT  1764 0 1764.56 4 ;
    END
  END wb_we_i
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER Metal4 ;
        RECT 97.805 45 100.305 2349.2 ;
        RECT 185.805 45 188.305 2349.2 ;
        RECT 273.805 45 276.305 2349.2 ;
        RECT 361.805 45 364.305 2349.2 ;
        RECT 449.805 45 452.305 2349.2 ;
        RECT 537.8050000000001 45 540.3050000000001 2349.2 ;
        RECT 625.8050000000001 45 628.3050000000001 2349.2 ;
        RECT 713.8050000000001 45 716.3050000000001 2349.2 ;
        RECT 801.8050000000001 45 804.3050000000001 2349.2 ;
        RECT 889.8050000000001 45 892.3050000000001 2349.2 ;
        RECT 977.8050000000001 45 980.3050000000001 2349.2 ;
        RECT 1065.805 45 1068.305 2349.2 ;
        RECT 1153.805 45 1156.305 2349.2 ;
        RECT 1241.805 45 1244.305 2349.2 ;
        RECT 1329.805 45 1332.305 2349.2 ;
        RECT 1417.805 45 1420.305 2349.2 ;
        RECT 1505.805 45 1508.305 2349.2 ;
        RECT 1593.805 45 1596.305 2349.2 ;
        RECT 1681.805 45 1684.305 2349.2 ;
        RECT 1769.805 45 1772.305 2349.2 ;
        RECT 1857.805 45 1860.305 2349.2 ;
        RECT 1945.805 45 1948.305 2349.2 ;
        RECT 2033.805 45 2036.305 2349.2 ;
        RECT 2121.805 45 2124.305 2349.2 ;

        RECT  2145.96 811.14 2147.56 1533.02 ;
        RECT  2044.6 1575.54 2046.2 2305.26 ;
        RECT  2145.96 42.82 2147.56 764.7 ;
        RECT  1956.68 1575.54 1958.28 2305.26 ;
        RECT  2044.6 38.9 2046.2 768.62 ;
        RECT  1956.68 807.22 1958.28 1536.94 ;
        RECT  2145.96 1579.46 2147.56 2301.34 ;
        RECT  2044.6 807.22 2046.2 1536.94 ;
        RECT  1956.68 38.9 1958.28 768.62 ;
        RECT  1868.2 38.9 1869.8 768.62 ;
        RECT  1780.28 807.22 1781.88 1536.94 ;
        RECT  1692.36 1575.54 1693.96 2305.26 ;
        RECT  1868.2 807.22 1869.8 1536.94 ;
        RECT  1780.28 38.9 1781.88 768.62 ;
        RECT  1604.44 1575.54 1606.04 2305.26 ;
        RECT  1868.2 1575.54 1869.8 2305.26 ;
        RECT  1692.36 38.9 1693.96 768.62 ;
        RECT  1604.44 807.22 1606.04 1536.94 ;
        RECT  1780.28 1575.54 1781.88 2305.26 ;
        RECT  1692.36 807.22 1693.96 1536.94 ;
        RECT  1604.44 38.9 1606.04 768.62 ;
        RECT  1516.52 38.9 1518.12 768.62 ;
        RECT  1428.6 807.22 1430.2 1536.94 ;
        RECT  1516.52 807.22 1518.12 1536.94 ;
        RECT  1428.6 38.9 1430.2 768.62 ;
        RECT  1252.2 1575.54 1253.8 2305.26 ;
        RECT  1516.52 1575.54 1518.12 2305.26 ;
        RECT  1252.2 807.22 1253.8 1536.94 ;
        RECT  1428.6 1575.54 1430.2 2305.26 ;
        RECT  1252.2 38.9 1253.8 768.62 ;
        RECT  1076.36 38.9 1077.96 768.62 ;
        RECT  993.48 811.14 995.08 1533.02 ;
        RECT  900.52 1575.54 902.12 2305.26 ;
        RECT  1076.36 807.22 1077.96 1536.94 ;
        RECT  993.48 42.82 995.08 764.7 ;
        RECT  812.6 1575.54 814.2 2305.26 ;
        RECT  1076.36 1575.54 1077.96 2305.26 ;
        RECT  900.52 38.9 902.12 768.62 ;
        RECT  812.6 807.22 814.2 1536.94 ;
        RECT  993.48 1579.46 995.08 2301.34 ;
        RECT  900.52 807.22 902.12 1536.94 ;
        RECT  812.6 38.9 814.2 768.62 ;
        RECT  724.68 38.9 726.28 768.62 ;
        RECT  636.2 807.22 637.8 1536.94 ;
        RECT  548.28 1575.54 549.88 2305.26 ;
        RECT  724.68 807.22 726.28 1536.94 ;
        RECT  636.2 38.9 637.8 768.62 ;
        RECT  460.36 1575.54 461.96 2305.26 ;
        RECT  724.68 1575.54 726.28 2305.26 ;
        RECT  548.28 38.9 549.88 768.62 ;
        RECT  460.36 807.22 461.96 1536.94 ;
        RECT  636.2 1575.54 637.8 2305.26 ;
        RECT  548.28 807.22 549.88 1536.94 ;
        RECT  460.36 38.9 461.96 768.62 ;
        RECT  372.44 38.9 374.04 768.62 ;
        RECT  284.52 807.22 286.12 1536.94 ;
        RECT  196.6 1575.54 198.2 2305.26 ;
        RECT  372.44 807.22 374.04 1536.94 ;
        RECT  284.52 38.9 286.12 768.62 ;
        RECT  108.68 1575.54 110.28 2305.26 ;
        RECT  372.44 1575.54 374.04 2305.26 ;
        RECT  196.6 38.9 198.2 768.62 ;
        RECT  108.68 807.22 110.28 1536.94 ;
        RECT  284.52 1575.54 286.12 2305.26 ;
        RECT  196.6 807.22 198.2 1536.94 ;
        RECT  108.68 38.9 110.28 768.62 ;
        RECT  2115.92 2298.515 2117.52 2352.3 ;
        RECT  2115.92 1530.515 2117.52 1580.44 ;
        RECT  2115.92 762.515 2117.52 812.44 ;
        RECT  2115.92 15.38 2117.52 44.44 ;
        RECT  1925.92 2298.49 1927.52 2352.3 ;
        RECT  1925.92 1530.49 1927.52 1585.075 ;
        RECT  1925.92 762.49 1927.52 817.075 ;
        RECT  1925.92 15.38 1927.52 49.075 ;
        RECT  1735.92 2298.49 1737.52 2352.3 ;
        RECT  1735.92 1530.49 1737.52 1585.075 ;
        RECT  1735.92 762.49 1737.52 817.075 ;
        RECT  1735.92 15.38 1737.52 49.075 ;
        RECT  1545.92 2298.515 1547.52 2352.3 ;
        RECT  1545.92 1530.515 1547.52 1580.44 ;
        RECT  1545.92 762.515 1547.52 812.44 ;
        RECT  1545.92 15.38 1547.52 44.44 ;
        RECT  1355.92 15.38 1357.52 2352.3 ;
        RECT  1165.92 15.38 1167.52 2352.3 ;
        RECT  975.92 15.38 977.52 44.44 ;
        RECT  785.92 2298.515 787.52 2352.3 ;
        RECT  785.92 1530.515 787.52 1585.075 ;
        RECT  785.92 762.515 787.52 817.075 ;
        RECT  785.92 15.38 787.52 49.075 ;
        RECT  595.92 2298.49 597.52 2352.3 ;
        RECT  595.92 1530.49 597.52 1585.075 ;
        RECT  595.92 762.49 597.52 817.075 ;
        RECT  595.92 15.38 597.52 49.075 ;
        RECT  405.92 2298.49 407.52 2352.3 ;
        RECT  405.92 1530.49 407.52 1585.05 ;
        RECT  405.92 762.49 407.52 817.05 ;
        RECT  405.92 15.38 407.52 49.05 ;
        RECT  215.92 15.38 217.52 44.44 ;
        RECT  25.92 15.38 27.52 2352.3 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER Metal4 ;
        RECT 93.83500000000001 45 96.33500000000001 725 ;
        RECT 93.83500000000001 813 96.33500000000001 1493 ;
        RECT 93.83500000000001 1581 96.33500000000001 2261 ;
        RECT 40.0 45 42.5 2349.2 ;
        RECT 181.835 45 184.335 725 ;
        RECT 181.835 813 184.335 1493 ;
        RECT 181.835 1581 184.335 2261 ;
        RECT 128.0 45 130.5 2349.2 ;
        RECT 269.835 45 272.335 725 ;
        RECT 269.835 813 272.335 1493 ;
        RECT 269.835 1581 272.335 2261 ;
        RECT 216.0 45 218.5 2349.2 ;
        RECT 357.835 45 360.335 725 ;
        RECT 357.835 813 360.335 1493 ;
        RECT 357.835 1581 360.335 2261 ;
        RECT 304.0 45 306.5 2349.2 ;
        RECT 445.835 45 448.335 725 ;
        RECT 445.835 813 448.335 1493 ;
        RECT 445.835 1581 448.335 2261 ;
        RECT 392.0 45 394.5 2349.2 ;
        RECT 533.835 45 536.335 725 ;
        RECT 533.835 813 536.335 1493 ;
        RECT 533.835 1581 536.335 2261 ;
        RECT 480.0 45 482.5 2349.2 ;
        RECT 621.835 45 624.335 725 ;
        RECT 621.835 813 624.335 1493 ;
        RECT 621.835 1581 624.335 2261 ;
        RECT 568.0 45 570.5 2349.2 ;
        RECT 709.835 45 712.335 725 ;
        RECT 709.835 813 712.335 1493 ;
        RECT 709.835 1581 712.335 2261 ;
        RECT 656.0 45 658.5 2349.2 ;
        RECT 797.835 45 800.335 725 ;
        RECT 797.835 813 800.335 1493 ;
        RECT 797.835 1581 800.335 2261 ;
        RECT 744.0 45 746.5 2349.2 ;
        RECT 885.835 45 888.335 725 ;
        RECT 885.835 813 888.335 1493 ;
        RECT 885.835 1581 888.335 2261 ;
        RECT 832.0 45 834.5 2349.2 ;
        RECT 973.835 45 976.335 725 ;
        RECT 973.835 813 976.335 1493 ;
        RECT 973.835 1581 976.335 2261 ;
        RECT 920.0 45 922.5 2349.2 ;
        RECT 1061.835 45 1064.335 725 ;
        RECT 1061.835 813 1064.335 1493 ;
        RECT 1061.835 1581 1064.335 2261 ;
        RECT 1008.0 45 1010.5 2349.2 ;
        RECT 1149.835 45 1152.335 725 ;
        RECT 1149.835 813 1152.335 1493 ;
        RECT 1149.835 1581 1152.335 2261 ;
        RECT 1096.0 45 1098.5 2349.2 ;
        RECT 1237.835 45 1240.335 725 ;
        RECT 1237.835 813 1240.335 1493 ;
        RECT 1237.835 1581 1240.335 2261 ;
        RECT 1184.0 45 1186.5 2349.2 ;
        RECT 1325.835 45 1328.335 725 ;
        RECT 1325.835 813 1328.335 1493 ;
        RECT 1325.835 1581 1328.335 2261 ;
        RECT 1272.0 45 1274.5 2349.2 ;
        RECT 1413.835 45 1416.335 725 ;
        RECT 1413.835 813 1416.335 1493 ;
        RECT 1413.835 1581 1416.335 2261 ;
        RECT 1360.0 45 1362.5 2349.2 ;
        RECT 1501.835 45 1504.335 725 ;
        RECT 1501.835 813 1504.335 1493 ;
        RECT 1501.835 1581 1504.335 2261 ;
        RECT 1448.0 45 1450.5 2349.2 ;
        RECT 1589.835 45 1592.335 725 ;
        RECT 1589.835 813 1592.335 1493 ;
        RECT 1589.835 1581 1592.335 2261 ;
        RECT 1536.0 45 1538.5 2349.2 ;
        RECT 1677.835 45 1680.335 725 ;
        RECT 1677.835 813 1680.335 1493 ;
        RECT 1677.835 1581 1680.335 2261 ;
        RECT 1624.0 45 1626.5 2349.2 ;
        RECT 1765.835 45 1768.335 725 ;
        RECT 1765.835 813 1768.335 1493 ;
        RECT 1765.835 1581 1768.335 2261 ;
        RECT 1712.0 45 1714.5 2349.2 ;
        RECT 1853.835 45 1856.335 725 ;
        RECT 1853.835 813 1856.335 1493 ;
        RECT 1853.835 1581 1856.335 2261 ;
        RECT 1800.0 45 1802.5 2349.2 ;
        RECT 1941.835 45 1944.335 725 ;
        RECT 1941.835 813 1944.335 1493 ;
        RECT 1941.835 1581 1944.335 2261 ;
        RECT 1888.0 45 1890.5 2349.2 ;
        RECT 2029.835 45 2032.335 725 ;
        RECT 2029.835 813 2032.335 1493 ;
        RECT 2029.835 1581 2032.335 2261 ;
        RECT 1976.0 45 1978.5 2349.2 ;
        RECT 2117.835 45 2120.335 725 ;
        RECT 2117.835 813 2120.335 1493 ;
        RECT 2117.835 1581 2120.335 2261 ;
        RECT 2064.0 45 2066.5 2349.2 ;

        RECT  2054.68 1575.54 2056.28 2305.26 ;
        RECT  1966.76 1575.54 1968.36 2305.26 ;
        RECT  2054.68 38.9 2056.28 768.62 ;
        RECT  1966.76 807.22 1968.36 1536.94 ;
        RECT  2054.68 807.22 2056.28 1536.94 ;
        RECT  1966.76 38.9 1968.36 768.62 ;
        RECT  1878.28 38.9 1879.88 768.62 ;
        RECT  1790.36 807.22 1791.96 1536.94 ;
        RECT  1702.44 1575.54 1704.04 2305.26 ;
        RECT  1878.28 807.22 1879.88 1536.94 ;
        RECT  1790.36 38.9 1791.96 768.62 ;
        RECT  1614.52 1575.54 1616.12 2305.26 ;
        RECT  1878.28 1575.54 1879.88 2305.26 ;
        RECT  1702.44 38.9 1704.04 768.62 ;
        RECT  1614.52 807.22 1616.12 1536.94 ;
        RECT  1790.36 1575.54 1791.96 2305.26 ;
        RECT  1702.44 807.22 1704.04 1536.94 ;
        RECT  1614.52 38.9 1616.12 768.62 ;
        RECT  1526.6 38.9 1528.2 768.62 ;
        RECT  1438.68 807.22 1440.28 1536.94 ;
        RECT  1345.16 1575.54 1346.76 2305.26 ;
        RECT  1526.6 807.22 1528.2 1536.94 ;
        RECT  1438.68 38.9 1440.28 768.62 ;
        RECT  1262.28 1575.54 1263.88 2305.26 ;
        RECT  1526.6 1575.54 1528.2 2305.26 ;
        RECT  1345.16 38.9 1346.76 768.62 ;
        RECT  1262.28 807.22 1263.88 1536.94 ;
        RECT  1438.68 1575.54 1440.28 2305.26 ;
        RECT  1345.16 807.22 1346.76 1536.94 ;
        RECT  1262.28 38.9 1263.88 768.62 ;
        RECT  1086.44 38.9 1088.04 768.62 ;
        RECT  910.6 1575.54 912.2 2305.26 ;
        RECT  1086.44 807.22 1088.04 1536.94 ;
        RECT  822.68 1575.54 824.28 2305.26 ;
        RECT  1086.44 1575.54 1088.04 2305.26 ;
        RECT  910.6 38.9 912.2 768.62 ;
        RECT  822.68 807.22 824.28 1536.94 ;
        RECT  910.6 807.22 912.2 1536.94 ;
        RECT  822.68 38.9 824.28 768.62 ;
        RECT  734.76 38.9 736.36 768.62 ;
        RECT  646.28 807.22 647.88 1536.94 ;
        RECT  558.36 1575.54 559.96 2305.26 ;
        RECT  734.76 807.22 736.36 1536.94 ;
        RECT  646.28 38.9 647.88 768.62 ;
        RECT  470.44 1575.54 472.04 2305.26 ;
        RECT  734.76 1575.54 736.36 2305.26 ;
        RECT  558.36 38.9 559.96 768.62 ;
        RECT  470.44 807.22 472.04 1536.94 ;
        RECT  646.28 1575.54 647.88 2305.26 ;
        RECT  558.36 807.22 559.96 1536.94 ;
        RECT  470.44 38.9 472.04 768.62 ;
        RECT  382.52 38.9 384.12 768.62 ;
        RECT  294.6 807.22 296.2 1536.94 ;
        RECT  206.68 1575.54 208.28 2305.26 ;
        RECT  382.52 807.22 384.12 1536.94 ;
        RECT  294.6 38.9 296.2 768.62 ;
        RECT  118.76 1575.54 120.36 2305.26 ;
        RECT  382.52 1575.54 384.12 2305.26 ;
        RECT  206.68 38.9 208.28 768.62 ;
        RECT  118.76 807.22 120.36 1536.94 ;
        RECT  294.6 1575.54 296.2 2305.26 ;
        RECT  206.68 807.22 208.28 1536.94 ;
        RECT  118.76 38.9 120.36 768.62 ;
        RECT  2125.52 15.38 2127.12 2352.3 ;
        RECT  1935.52 2298.515 1937.12 2352.3 ;
        RECT  1935.52 1530.515 1937.12 1585.075 ;
        RECT  1935.52 762.515 1937.12 817.075 ;
        RECT  1935.52 15.38 1937.12 49.075 ;
        RECT  1745.52 2298.49 1747.12 2352.3 ;
        RECT  1745.52 1530.49 1747.12 1585.075 ;
        RECT  1745.52 762.49 1747.12 817.075 ;
        RECT  1745.52 15.38 1747.12 49.075 ;
        RECT  1555.52 2298.49 1557.12 2352.3 ;
        RECT  1555.52 1530.49 1557.12 1585.075 ;
        RECT  1555.52 762.49 1557.12 817.075 ;
        RECT  1555.52 15.38 1557.12 49.075 ;
        RECT  1365.52 2298.515 1367.12 2352.3 ;
        RECT  1365.52 1530.515 1367.12 1580.44 ;
        RECT  1365.52 762.515 1367.12 812.44 ;
        RECT  1365.52 15.38 1367.12 44.44 ;
        RECT  1175.52 15.38 1177.12 2352.3 ;
        RECT  985.52 15.38 987.12 2352.3 ;
        RECT  795.52 2298.515 797.12 2352.3 ;
        RECT  795.52 1530.515 797.12 1585.05 ;
        RECT  795.52 762.515 797.12 817.05 ;
        RECT  795.52 15.38 797.12 49.05 ;
        RECT  605.52 2298.49 607.12 2352.3 ;
        RECT  605.52 1530.49 607.12 1585.075 ;
        RECT  605.52 762.49 607.12 817.075 ;
        RECT  605.52 15.38 607.12 49.075 ;
        RECT  415.52 2298.49 417.12 2352.3 ;
        RECT  415.52 1530.49 417.12 1585.075 ;
        RECT  415.52 762.49 417.12 817.075 ;
        RECT  415.52 15.38 417.12 49.075 ;
        RECT  225.52 2298.515 227.12 2352.3 ;
        RECT  225.52 1530.515 227.12 1580.44 ;
        RECT  225.52 762.515 227.12 812.44 ;
        RECT  225.52 15.38 227.12 44.44 ;
        RECT  35.52 15.38 37.12 2352.3 ;
    END
  END VSS
  OBS
    LAYER Pwell ;
     RECT  0 0 2175 2352.3 ;
    LAYER Nwell ;
     RECT  0 0 2175 2352.3 ;
    LAYER Metal1 ;
     RECT  0 0 2175 2352.3 ;
    LAYER Metal2 ;
     RECT  0 0 2175 2352.3 ;
    LAYER Metal3 ;
     RECT  0 0 2175 2352.3 ;
    LAYER Metal4 ;
     RECT  0 0 2175 2352.3 ;
    LAYER Metal5 ;
        RECT 10 0 2165 34.5 ;
        RECT 10 49.5 2165 79.5 ;
        RECT 10 94.5 2165 124.5 ;
        RECT 10 139.5 2165 169.5 ;
        RECT 10 184.5 2165 214.5 ;
        RECT 10 229.5 2165 259.5 ;
        RECT 10 274.5 2165 304.5 ;
        RECT 10 319.5 2165 349.5 ;
        RECT 10 364.5 2165 394.5 ;
        RECT 10 409.5 2165 439.5 ;
        RECT 10 454.5 2165 484.5 ;
        RECT 10 499.5 2165 529.5 ;
        RECT 10 544.5 2165 574.5 ;
        RECT 10 589.5 2165 619.5 ;
        RECT 10 634.5 2165 664.5 ;
        RECT 10 679.5 2165 709.5 ;
        RECT 10 724.5 2165 754.5 ;
        RECT 10 769.5 2165 799.5 ;
        RECT 10 814.5 2165 844.5 ;
        RECT 10 859.5 2165 889.5 ;
        RECT 10 904.5 2165 934.5 ;
        RECT 10 949.5 2165 979.5 ;
        RECT 10 994.5 2165 1024.5 ;
        RECT 10 1039.5 2165 1069.5 ;
        RECT 10 1084.5 2165 1114.5 ;
        RECT 10 1129.5 2165 1159.5 ;
        RECT 10 1174.5 2165 1204.5 ;
        RECT 10 1219.5 2165 1249.5 ;
        RECT 10 1264.5 2165 1294.5 ;
        RECT 10 1309.5 2165 1339.5 ;
        RECT 10 1354.5 2165 1384.5 ;
        RECT 10 1399.5 2165 1429.5 ;
        RECT 10 1444.5 2165 1474.5 ;
        RECT 10 1489.5 2165 1519.5 ;
        RECT 10 1534.5 2165 1564.5 ;
        RECT 10 1579.5 2165 1609.5 ;
        RECT 10 1624.5 2165 1654.5 ;
        RECT 10 1669.5 2165 1699.5 ;
        RECT 10 1714.5 2165 1744.5 ;
        RECT 10 1759.5 2165 1789.5 ;
        RECT 10 1804.5 2165 1834.5 ;
        RECT 10 1849.5 2165 1879.5 ;
        RECT 10 1894.5 2165 1924.5 ;
        RECT 10 1939.5 2165 1969.5 ;
        RECT 10 1984.5 2165 2014.5 ;
        RECT 10 2029.5 2165 2059.5 ;
        RECT 10 2074.5 2165 2104.5 ;
        RECT 10 2119.5 2165 2149.5 ;
        RECT 10 2164.5 2165 2194.5 ;
        RECT 10 2209.5 2165 2239.5 ;
        RECT 10 2254.5 2165 2284.5 ;
        RECT 10 2299.5 2165 2329.5 ;
  END
END efuse_ctrl
END LIBRARY
