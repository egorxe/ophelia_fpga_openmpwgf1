.subckt efuse_bitcell  select anode VSS
X0 anode net1 efuse
X1 net1 select VSS VSS nfet_06v0 L=0.70u W=50u
.ends

.subckt efuse_bitcell2  select anode VSS
X0 net1 anode efuse
X1 net1 select VSS VSS nfet_06v0 L=0.70u W=50u
.ends

.subckt efuse_sense_amp  VDD nPRESET OUT SENSE VSS FUSE
X2 net1 nPRESET VDD VDD pfet_06v0 L=0.50u W=1.9u
x1 net2 OUT VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__inv_2
x2 net1 net2 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__inv_1
x3 net2 net1 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__inv_1
X1 net1 SENSE FUSE VSS nfet_06v0 L=0.60u W=0.5u
.ends

.subckt efuse_byte ANODE_0 ANODE_1 ANODE_2 ANODE_3 ANODE_4 ANODE_5 ANODE_6 ANODE_7 VSS LINE_SEL
x0 LINE_SEL ANODE_0 VSS efuse_bitcell2
x1 LINE_SEL ANODE_1 VSS efuse_bitcell
x2 LINE_SEL ANODE_2 VSS efuse_bitcell
x3 LINE_SEL ANODE_3 VSS efuse_bitcell2
x4 LINE_SEL ANODE_4 VSS efuse_bitcell2
x5 LINE_SEL ANODE_5 VSS efuse_bitcell
x6 LINE_SEL ANODE_6 VSS efuse_bitcell
x7 LINE_SEL ANODE_7 VSS efuse_bitcell2
.ends

.subckt efuse_array LINE[0] LINE[1] LINE[2] LINE[3] LINE[4] LINE[5] LINE[6] LINE[7] LINE[8] LINE[9] LINE[10] LINE[11] LINE[12] LINE[13] LINE[14] LINE[15] VDD VSS COL_PROG[0] COL_PROG[1] COL_PROG[2] COL_PROG[3] COL_PROG[4] COL_PROG[5] COL_PROG[6] COL_PROG[7] SENSE nPRESET DO[0] DO[1] DO[2] DO[3] DO[4] DO[5] DO[6] DO[7] 
x0_0 net0 net1 net2 net3 net4 net5 net6 net7 VSS LINE_0_buf efuse_byte
x4_0 LINE[0] LINE_0_buf VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__buf_1
x0_1 net0 net1 net2 net3 net4 net5 net6 net7 VSS LINE_1_buf efuse_byte
x4_1 LINE[1] LINE_1_buf VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__buf_1
x0_2 net0 net1 net2 net3 net4 net5 net6 net7 VSS LINE_2_buf efuse_byte
x4_2 LINE[2] LINE_2_buf VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__buf_1
x0_3 net0 net1 net2 net3 net4 net5 net6 net7 VSS LINE_3_buf efuse_byte
x4_3 LINE[3] LINE_3_buf VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__buf_1
x0_4 net0 net1 net2 net3 net4 net5 net6 net7 VSS LINE_4_buf efuse_byte
x4_4 LINE[4] LINE_4_buf VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__buf_1
x0_5 net0 net1 net2 net3 net4 net5 net6 net7 VSS LINE_5_buf efuse_byte
x4_5 LINE[5] LINE_5_buf VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__buf_1
x0_6 net0 net1 net2 net3 net4 net5 net6 net7 VSS LINE_6_buf efuse_byte
x4_6 LINE[6] LINE_6_buf VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__buf_1
x0_7 net0 net1 net2 net3 net4 net5 net6 net7 VSS LINE_7_buf efuse_byte
x4_7 LINE[7] LINE_7_buf VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__buf_1
x0_8 net0 net1 net2 net3 net4 net5 net6 net7 VSS LINE_8_buf efuse_byte
x4_8 LINE[8] LINE_8_buf VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__buf_1
x0_9 net0 net1 net2 net3 net4 net5 net6 net7 VSS LINE_9_buf efuse_byte
x4_9 LINE[9] LINE_9_buf VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__buf_1
x0_10 net0 net1 net2 net3 net4 net5 net6 net7 VSS LINE_10_buf efuse_byte
x4_10 LINE[10] LINE_10_buf VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__buf_1
x0_11 net0 net1 net2 net3 net4 net5 net6 net7 VSS LINE_11_buf efuse_byte
x4_11 LINE[11] LINE_11_buf VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__buf_1
x0_12 net0 net1 net2 net3 net4 net5 net6 net7 VSS LINE_12_buf efuse_byte
x4_12 LINE[12] LINE_12_buf VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__buf_1
x0_13 net0 net1 net2 net3 net4 net5 net6 net7 VSS LINE_13_buf efuse_byte
x4_13 LINE[13] LINE_13_buf VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__buf_1
x0_14 net0 net1 net2 net3 net4 net5 net6 net7 VSS LINE_14_buf efuse_byte
x4_14 LINE[14] LINE_14_buf VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__buf_1
x0_15 net0 net1 net2 net3 net4 net5 net6 net7 VSS LINE_15_buf efuse_byte
x4_15 LINE[15] LINE_15_buf VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__buf_1

X0 net0 COL_PROG[0] VDD VDD pfet_06v0 L=0.50u W=50u

X1 net1 COL_PROG[1] VDD VDD pfet_06v0 L=0.50u W=50u

X2 net2 COL_PROG[2] VDD VDD pfet_06v0 L=0.50u W=50u

X3 net3 COL_PROG[3] VDD VDD pfet_06v0 L=0.50u W=50u

X4 net4 COL_PROG[4] VDD VDD pfet_06v0 L=0.50u W=50u

X5 net5 COL_PROG[5] VDD VDD pfet_06v0 L=0.50u W=50u

X6 net6 COL_PROG[6] VDD VDD pfet_06v0 L=0.50u W=50u

X7 net7 COL_PROG[7] VDD VDD pfet_06v0 L=0.50u W=50u

x1_0 VDD nPRESET DO_0_buf SENSE VSS net0 efuse_sense_amp
x3_0 DO_0_buf DO[0] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__buf_1
x1_1 VDD nPRESET DO_1_buf SENSE VSS net1 efuse_sense_amp
x3_1 DO_1_buf DO[1] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__buf_1
x1_2 VDD nPRESET DO_2_buf SENSE VSS net2 efuse_sense_amp
x3_2 DO_2_buf DO[2] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__buf_1
x1_3 VDD nPRESET DO_3_buf SENSE VSS net3 efuse_sense_amp
x3_3 DO_3_buf DO[3] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__buf_1
x1_4 VDD nPRESET DO_4_buf SENSE VSS net4 efuse_sense_amp
x3_4 DO_4_buf DO[4] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__buf_1
x1_5 VDD nPRESET DO_5_buf SENSE VSS net5 efuse_sense_amp
x3_5 DO_5_buf DO[5] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__buf_1
x1_6 VDD nPRESET DO_6_buf SENSE VSS net6 efuse_sense_amp
x3_6 DO_6_buf DO[6] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__buf_1
x1_7 VDD nPRESET DO_7_buf SENSE VSS net7 efuse_sense_amp
x3_7 DO_7_buf DO[7] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__buf_1
x2_0 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
x2_1 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
x2_2 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
x2_3 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
x2_4 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
x2_5 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
x2_6 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
x2_7 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
x2_8 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
x2_9 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
x2_10 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
x2_11 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
x2_12 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
x2_13 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
x2_14 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
x2_15 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
x2_16 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
x2_17 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
x2_18 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
x2_19 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
x2_20 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
x2_21 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
x2_22 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
x2_23 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
x2_24 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
x2_25 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
x2_26 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
x2_27 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
x2_28 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
x2_29 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
x2_30 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
x2_31 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
x2_32 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
x2_33 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
x2_34 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
x2_35 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
x2_36 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
x2_37 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
x2_38 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
x2_39 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
x2_40 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
x2_41 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
x2_42 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
x2_43 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
x2_44 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
x2_45 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
x2_46 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
x2_47 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
x2_48 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
x2_49 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
x2_50 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
x2_51 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
x2_52 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
x2_53 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
x2_54 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
x2_55 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
x2_56 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
x2_57 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
x2_58 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
x2_59 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
x2_60 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
x2_61 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
x2_62 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
x2_63 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
x2_64 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
x2_65 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
x2_66 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
x2_67 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
x2_68 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
x2_69 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
x2_70 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
x2_71 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
x2_72 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
x2_73 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
x2_74 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
x2_75 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
x2_76 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
x2_77 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
x2_78 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
x2_79 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
x2_80 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
x2_81 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
x2_82 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
x2_83 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
x2_84 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
x2_85 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
x2_86 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
x2_87 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
x2_88 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
x2_89 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
x2_90 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
x2_91 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
x2_92 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
x2_93 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
x2_94 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
x2_95 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
x2_96 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
x2_97 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
x2_98 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
x2_99 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
x2_100 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
x2_101 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
x2_102 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
x2_103 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
x2_104 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
x2_105 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
x2_106 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
x2_107 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
x2_108 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
x2_109 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
x2_110 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
x2_111 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
x2_112 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
x2_113 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
x2_114 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
x2_115 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
x2_116 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
x2_117 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
x2_118 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
x2_119 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
x2_120 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
x2_121 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
x2_122 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
x2_123 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
x2_124 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
x2_125 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
x2_126 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
x2_127 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
x2_128 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
x2_129 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
x2_130 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
x2_131 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
x2_132 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
x2_133 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
x2_134 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
x2_135 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
x2_136 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
x2_137 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
x2_138 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
x2_139 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
x2_140 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
x2_141 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
x2_142 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
x2_143 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
x2_144 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
x2_145 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
x2_146 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
x2_147 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
x2_148 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
x2_149 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
x2_150 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
x2_151 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
x2_152 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
x2_153 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
x2_154 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
x2_155 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
x2_156 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
x2_157 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
x2_158 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
x2_159 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
x2_160 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
x2_161 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
x2_162 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
x2_163 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
x2_164 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
x2_165 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
x2_166 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
x2_167 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
x2_168 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
x2_169 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
x2_170 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
x2_171 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
x2_172 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
x2_173 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
x2_174 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
x2_175 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
x2_176 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
x2_177 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
x2_178 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
x2_179 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
x2_180 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
x2_181 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
x2_182 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
x2_183 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
x2_184 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
x2_185 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
x2_186 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
x2_187 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
x2_188 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
x2_189 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
x2_190 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
x2_191 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
x2_192 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
x2_193 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
x2_194 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
x2_195 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
x2_196 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
x2_197 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
x2_198 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
x2_199 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
x2_200 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
x2_201 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
x2_202 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
x2_203 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
x2_204 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
x2_205 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
x2_206 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
x2_207 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
x2_208 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
x2_209 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
.ends

.end
