VERSION 5.8 ;
BUSBITCHARS "[]" ;
DIVIDERCHAR "/" ;
UNITS
    DATABASE MICRONS 2000 ;
END UNITS
MACRO efuse_ctrl
  FOREIGN efuse_ctrl 0 0 ;
  CLASS BLOCK ;
  ORIGIN 0 0 ;
  SIZE 2175 BY 2352.3 ;
  PIN wb_ack_o
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT  1884.96 0 1885.52 4 ;
    END
  END wb_ack_o
  PIN wb_adr_i[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT  33.6 0 34.16 4 ;
    END
  END wb_adr_i[0]
  PIN wb_adr_i[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT  672 0 672.56 4 ;
    END
  END wb_adr_i[10]
  PIN wb_adr_i[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT  97.44 0 98 4 ;
    END
  END wb_adr_i[1]
  PIN wb_adr_i[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT  161.28 0 161.84 4 ;
    END
  END wb_adr_i[2]
  PIN wb_adr_i[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT  225.12 0 225.68 4 ;
    END
  END wb_adr_i[3]
  PIN wb_adr_i[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT  288.96 0 289.52 4 ;
    END
  END wb_adr_i[4]
  PIN wb_adr_i[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT  352.8 0 353.36 4 ;
    END
  END wb_adr_i[5]
  PIN wb_adr_i[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT  416.64 0 417.2 4 ;
    END
  END wb_adr_i[6]
  PIN wb_adr_i[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT  480.48 0 481.04 4 ;
    END
  END wb_adr_i[7]
  PIN wb_adr_i[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT  544.32 0 544.88 4 ;
    END
  END wb_adr_i[8]
  PIN wb_adr_i[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT  608.16 0 608.72 4 ;
    END
  END wb_adr_i[9]
  PIN wb_clk_i
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT  2076.48 0 2077.04 4 ;
    END
  END wb_clk_i
  PIN wb_cyc_i
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT  2012.64 0 2013.2 4 ;
    END
  END wb_cyc_i
  PIN wb_dat_i[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT  1246.56 0 1247.12 4 ;
    END
  END wb_dat_i[0]
  PIN wb_dat_i[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT  1310.4 0 1310.96 4 ;
    END
  END wb_dat_i[1]
  PIN wb_dat_i[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT  1374.24 0 1374.8 4 ;
    END
  END wb_dat_i[2]
  PIN wb_dat_i[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT  1438.08 0 1438.64 4 ;
    END
  END wb_dat_i[3]
  PIN wb_dat_i[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT  1501.92 0 1502.48 4 ;
    END
  END wb_dat_i[4]
  PIN wb_dat_i[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT  1565.76 0 1566.32 4 ;
    END
  END wb_dat_i[5]
  PIN wb_dat_i[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT  1629.6 0 1630.16 4 ;
    END
  END wb_dat_i[6]
  PIN wb_dat_i[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT  1693.44 0 1694 4 ;
    END
  END wb_dat_i[7]
  PIN wb_dat_o[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT  735.84 0 736.4 4 ;
    END
  END wb_dat_o[0]
  PIN wb_dat_o[1]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT  799.68 0 800.24 4 ;
    END
  END wb_dat_o[1]
  PIN wb_dat_o[2]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT  863.52 0 864.08 4 ;
    END
  END wb_dat_o[2]
  PIN wb_dat_o[3]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT  927.36 0 927.92 4 ;
    END
  END wb_dat_o[3]
  PIN wb_dat_o[4]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT  991.2 0 991.76 4 ;
    END
  END wb_dat_o[4]
  PIN wb_dat_o[5]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT  1055.04 0 1055.6 4 ;
    END
  END wb_dat_o[5]
  PIN wb_dat_o[6]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT  1118.88 0 1119.44 4 ;
    END
  END wb_dat_o[6]
  PIN wb_dat_o[7]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT  1182.72 0 1183.28 4 ;
    END
  END wb_dat_o[7]
  PIN wb_rst_i
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT  2140.32 0 2140.88 4 ;
    END
  END wb_rst_i
  PIN wb_sel_i
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT  1948.8 0 1949.36 4 ;
    END
  END wb_sel_i
  PIN wb_stb_i
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT  1821.12 0 1821.68 4 ;
    END
  END wb_stb_i
  PIN wb_we_i
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT  1757.28 0 1757.84 4 ;
    END
  END wb_we_i
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER Metal4 ;
        RECT 101.5 45 104.0 2349.2 ;
        RECT 189.5 45 192.0 2349.2 ;
        RECT 277.5 45 280.0 2349.2 ;
        RECT 365.5 45 368.0 2349.2 ;
        RECT 453.5 45 456.0 2349.2 ;
        RECT 541.5 45 544.0 2349.2 ;
        RECT 629.5 45 632.0 2349.2 ;
        RECT 717.5 45 720.0 2349.2 ;
        RECT 805.5 45 808.0 2349.2 ;
        RECT 893.5 45 896.0 2349.2 ;
        RECT 981.5 45 984.0 2349.2 ;
        RECT 1069.5 45 1072.0 2349.2 ;
        RECT 1157.5 45 1160.0 2349.2 ;
        RECT 1245.5 45 1248.0 2349.2 ;
        RECT 1333.5 45 1336.0 2349.2 ;
        RECT 1421.5 45 1424.0 2349.2 ;
        RECT 1509.5 45 1512.0 2349.2 ;
        RECT 1597.5 45 1600.0 2349.2 ;
        RECT 1685.5 45 1688.0 2349.2 ;
        RECT 1773.5 45 1776.0 2349.2 ;
        RECT 1861.5 45 1864.0 2349.2 ;
        RECT 1949.5 45 1952.0 2349.2 ;
        RECT 2037.5 45 2040.0 2349.2 ;
        RECT 2125.5 45 2128.0 2349.2 ;

        RECT  2142.6 807.22 2144.2 1536.94 ;
        RECT  2046.28 1575.54 2047.88 2305.26 ;
        RECT  2142.6 38.9 2144.2 768.62 ;
        RECT  1958.36 1575.54 1959.96 2305.26 ;
        RECT  2046.28 38.9 2047.88 768.62 ;
        RECT  1958.36 807.22 1959.96 1536.94 ;
        RECT  2142.6 1575.54 2144.2 2305.26 ;
        RECT  2046.28 807.22 2047.88 1536.94 ;
        RECT  1958.36 38.9 1959.96 768.62 ;
        RECT  1870.44 38.9 1872.04 768.62 ;
        RECT  1782.52 807.22 1784.12 1536.94 ;
        RECT  1694.6 1575.54 1696.2 2305.26 ;
        RECT  1870.44 807.22 1872.04 1536.94 ;
        RECT  1782.52 38.9 1784.12 768.62 ;
        RECT  1606.12 1575.54 1607.72 2305.26 ;
        RECT  1870.44 1575.54 1872.04 2305.26 ;
        RECT  1694.6 38.9 1696.2 768.62 ;
        RECT  1606.12 807.22 1607.72 1536.94 ;
        RECT  1782.52 1575.54 1784.12 2305.26 ;
        RECT  1694.6 807.22 1696.2 1536.94 ;
        RECT  1606.12 38.9 1607.72 768.62 ;
        RECT  1518.2 38.9 1519.8 768.62 ;
        RECT  1430.28 807.22 1431.88 1536.94 ;
        RECT  1518.2 807.22 1519.8 1536.94 ;
        RECT  1430.28 38.9 1431.88 768.62 ;
        RECT  1254.44 1575.54 1256.04 2305.26 ;
        RECT  1518.2 1575.54 1519.8 2305.26 ;
        RECT  1254.44 807.22 1256.04 1536.94 ;
        RECT  1430.28 1575.54 1431.88 2305.26 ;
        RECT  1254.44 38.9 1256.04 768.62 ;
        RECT  1078.6 38.9 1080.2 768.62 ;
        RECT  995.16 811.14 996.76 1533.02 ;
        RECT  902.2 1575.54 903.8 2305.26 ;
        RECT  1078.6 807.22 1080.2 1536.94 ;
        RECT  995.16 42.82 996.76 764.7 ;
        RECT  814.28 1575.54 815.88 2305.26 ;
        RECT  1078.6 1575.54 1080.2 2305.26 ;
        RECT  902.2 38.9 903.8 768.62 ;
        RECT  814.28 807.22 815.88 1536.94 ;
        RECT  995.16 1579.46 996.76 2301.34 ;
        RECT  902.2 807.22 903.8 1536.94 ;
        RECT  814.28 38.9 815.88 768.62 ;
        RECT  726.36 38.9 727.96 768.62 ;
        RECT  638.44 807.22 640.04 1536.94 ;
        RECT  550.52 1575.54 552.12 2305.26 ;
        RECT  726.36 807.22 727.96 1536.94 ;
        RECT  638.44 38.9 640.04 768.62 ;
        RECT  462.6 1575.54 464.2 2305.26 ;
        RECT  726.36 1575.54 727.96 2305.26 ;
        RECT  550.52 38.9 552.12 768.62 ;
        RECT  462.6 807.22 464.2 1536.94 ;
        RECT  638.44 1575.54 640.04 2305.26 ;
        RECT  550.52 807.22 552.12 1536.94 ;
        RECT  462.6 38.9 464.2 768.62 ;
        RECT  374.12 38.9 375.72 768.62 ;
        RECT  286.2 807.22 287.8 1536.94 ;
        RECT  198.28 1575.54 199.88 2305.26 ;
        RECT  374.12 807.22 375.72 1536.94 ;
        RECT  286.2 38.9 287.8 768.62 ;
        RECT  110.36 1575.54 111.96 2305.26 ;
        RECT  374.12 1575.54 375.72 2305.26 ;
        RECT  198.28 38.9 199.88 768.62 ;
        RECT  110.36 807.22 111.96 1536.94 ;
        RECT  286.2 1575.54 287.8 2305.26 ;
        RECT  198.28 807.22 199.88 1536.94 ;
        RECT  110.36 38.9 111.96 768.62 ;
        RECT  2115.92 2299.53 2117.52 2352.3 ;
        RECT  2115.92 1531.53 2117.52 1582.27 ;
        RECT  2115.92 763.53 2117.52 814.27 ;
        RECT  2115.92 15.38 2117.52 46.27 ;
        RECT  1925.92 2299.51 1927.52 2352.3 ;
        RECT  1925.92 1531.51 1927.52 1582.27 ;
        RECT  1925.92 763.505 1927.52 814.27 ;
        RECT  1925.92 15.38 1927.52 46.27 ;
        RECT  1735.92 2299.51 1737.52 2352.3 ;
        RECT  1735.92 1531.51 1737.52 1582.27 ;
        RECT  1735.92 763.505 1737.52 814.27 ;
        RECT  1735.92 15.38 1737.52 46.27 ;
        RECT  1545.92 2299.53 1547.52 2352.3 ;
        RECT  1545.92 1531.53 1547.52 1580.04 ;
        RECT  1545.92 763.53 1547.52 811.72 ;
        RECT  1545.92 15.38 1547.52 43.72 ;
        RECT  1355.92 15.38 1357.52 2352.3 ;
        RECT  1165.92 15.38 1167.52 2352.3 ;
        RECT  975.92 2299.51 977.52 2352.3 ;
        RECT  975.92 1531.51 977.52 1582.25 ;
        RECT  975.92 763.505 977.52 814.245 ;
        RECT  975.92 15.38 977.52 46.245 ;
        RECT  785.92 2299.53 787.52 2352.3 ;
        RECT  785.92 1531.53 787.52 1582.27 ;
        RECT  785.92 763.53 787.52 814.27 ;
        RECT  785.92 15.38 787.52 46.27 ;
        RECT  595.92 2299.51 597.52 2352.3 ;
        RECT  595.92 1531.51 597.52 1582.27 ;
        RECT  595.92 763.505 597.52 814.27 ;
        RECT  595.92 15.38 597.52 46.27 ;
        RECT  405.92 2299.51 407.52 2352.3 ;
        RECT  405.92 1531.51 407.52 1582.25 ;
        RECT  405.92 763.505 407.52 814.245 ;
        RECT  405.92 15.38 407.52 46.245 ;
        RECT  215.92 15.38 217.52 43.72 ;
        RECT  25.92 15.38 27.52 2352.3 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER Metal4 ;
        RECT 40.0 45 42.5 2349.2 ;
        RECT 128.0 45 130.5 2349.2 ;
        RECT 216.0 45 218.5 2349.2 ;
        RECT 304.0 45 306.5 2349.2 ;
        RECT 392.0 45 394.5 2349.2 ;
        RECT 480.0 45 482.5 2349.2 ;
        RECT 568.0 45 570.5 2349.2 ;
        RECT 656.0 45 658.5 2349.2 ;
        RECT 744.0 45 746.5 2349.2 ;
        RECT 832.0 45 834.5 2349.2 ;
        RECT 920.0 45 922.5 2349.2 ;
        RECT 1008.0 45 1010.5 2349.2 ;
        RECT 1096.0 45 1098.5 2349.2 ;
        RECT 1184.0 45 1186.5 2349.2 ;
        RECT 1272.0 45 1274.5 2349.2 ;
        RECT 1360.0 45 1362.5 2349.2 ;
        RECT 1448.0 45 1450.5 2349.2 ;
        RECT 1536.0 45 1538.5 2349.2 ;
        RECT 1624.0 45 1626.5 2349.2 ;
        RECT 1712.0 45 1714.5 2349.2 ;
        RECT 1800.0 45 1802.5 2349.2 ;
        RECT 1888.0 45 1890.5 2349.2 ;
        RECT 1976.0 45 1978.5 2349.2 ;
        RECT 2064.0 45 2066.5 2349.2 ;

        RECT  2152.68 807.22 2154.28 1536.94 ;
        RECT  2056.36 1575.54 2057.96 2305.26 ;
        RECT  2152.68 38.9 2154.28 768.62 ;
        RECT  1968.44 1575.54 1970.04 2305.26 ;
        RECT  2056.36 38.9 2057.96 768.62 ;
        RECT  1968.44 807.22 1970.04 1536.94 ;
        RECT  2152.68 1575.54 2154.28 2305.26 ;
        RECT  2056.36 807.22 2057.96 1536.94 ;
        RECT  1968.44 38.9 1970.04 768.62 ;
        RECT  1880.52 38.9 1882.12 768.62 ;
        RECT  1792.6 807.22 1794.2 1536.94 ;
        RECT  1704.68 1575.54 1706.28 2305.26 ;
        RECT  1880.52 807.22 1882.12 1536.94 ;
        RECT  1792.6 38.9 1794.2 768.62 ;
        RECT  1616.2 1575.54 1617.8 2305.26 ;
        RECT  1880.52 1575.54 1882.12 2305.26 ;
        RECT  1704.68 38.9 1706.28 768.62 ;
        RECT  1616.2 807.22 1617.8 1536.94 ;
        RECT  1792.6 1575.54 1794.2 2305.26 ;
        RECT  1704.68 807.22 1706.28 1536.94 ;
        RECT  1616.2 38.9 1617.8 768.62 ;
        RECT  1528.28 38.9 1529.88 768.62 ;
        RECT  1440.36 807.22 1441.96 1536.94 ;
        RECT  1346.84 1575.54 1348.44 2305.26 ;
        RECT  1528.28 807.22 1529.88 1536.94 ;
        RECT  1440.36 38.9 1441.96 768.62 ;
        RECT  1264.52 1575.54 1266.12 2305.26 ;
        RECT  1528.28 1575.54 1529.88 2305.26 ;
        RECT  1346.84 38.9 1348.44 768.62 ;
        RECT  1264.52 807.22 1266.12 1536.94 ;
        RECT  1440.36 1575.54 1441.96 2305.26 ;
        RECT  1346.84 807.22 1348.44 1536.94 ;
        RECT  1264.52 38.9 1266.12 768.62 ;
        RECT  1088.68 38.9 1090.28 768.62 ;
        RECT  912.28 1575.54 913.88 2305.26 ;
        RECT  1088.68 807.22 1090.28 1536.94 ;
        RECT  824.36 1575.54 825.96 2305.26 ;
        RECT  1088.68 1575.54 1090.28 2305.26 ;
        RECT  912.28 38.9 913.88 768.62 ;
        RECT  824.36 807.22 825.96 1536.94 ;
        RECT  912.28 807.22 913.88 1536.94 ;
        RECT  824.36 38.9 825.96 768.62 ;
        RECT  736.44 38.9 738.04 768.62 ;
        RECT  648.52 807.22 650.12 1536.94 ;
        RECT  560.6 1575.54 562.2 2305.26 ;
        RECT  736.44 807.22 738.04 1536.94 ;
        RECT  648.52 38.9 650.12 768.62 ;
        RECT  472.68 1575.54 474.28 2305.26 ;
        RECT  736.44 1575.54 738.04 2305.26 ;
        RECT  560.6 38.9 562.2 768.62 ;
        RECT  472.68 807.22 474.28 1536.94 ;
        RECT  648.52 1575.54 650.12 2305.26 ;
        RECT  560.6 807.22 562.2 1536.94 ;
        RECT  472.68 38.9 474.28 768.62 ;
        RECT  384.2 38.9 385.8 768.62 ;
        RECT  296.28 807.22 297.88 1536.94 ;
        RECT  208.36 1575.54 209.96 2305.26 ;
        RECT  384.2 807.22 385.8 1536.94 ;
        RECT  296.28 38.9 297.88 768.62 ;
        RECT  120.44 1575.54 122.04 2305.26 ;
        RECT  384.2 1575.54 385.8 2305.26 ;
        RECT  208.36 38.9 209.96 768.62 ;
        RECT  120.44 807.22 122.04 1536.94 ;
        RECT  296.28 1575.54 297.88 2305.26 ;
        RECT  208.36 807.22 209.96 1536.94 ;
        RECT  120.44 38.9 122.04 768.62 ;
        RECT  2125.52 15.38 2127.12 43.72 ;
        RECT  1935.52 2299.53 1937.12 2352.3 ;
        RECT  1935.52 1531.53 1937.12 1582.27 ;
        RECT  1935.52 763.53 1937.12 814.27 ;
        RECT  1935.52 15.38 1937.12 46.27 ;
        RECT  1745.52 2299.51 1747.12 2352.3 ;
        RECT  1745.52 1531.51 1747.12 1582.27 ;
        RECT  1745.52 763.505 1747.12 814.27 ;
        RECT  1745.52 15.38 1747.12 46.27 ;
        RECT  1555.52 2299.51 1557.12 2352.3 ;
        RECT  1555.52 1531.51 1557.12 1582.27 ;
        RECT  1555.52 763.505 1557.12 814.27 ;
        RECT  1555.52 15.38 1557.12 46.27 ;
        RECT  1365.52 2299.53 1367.12 2352.3 ;
        RECT  1365.52 1531.53 1367.12 1579.72 ;
        RECT  1365.52 763.53 1367.12 811.72 ;
        RECT  1365.52 15.38 1367.12 43.72 ;
        RECT  1175.52 15.38 1177.12 2352.3 ;
        RECT  985.52 15.38 987.12 2352.3 ;
        RECT  795.52 2299.53 797.12 2352.3 ;
        RECT  795.52 1531.53 797.12 1582.27 ;
        RECT  795.52 763.53 797.12 814.27 ;
        RECT  795.52 15.38 797.12 46.27 ;
        RECT  605.52 2299.51 607.12 2352.3 ;
        RECT  605.52 1531.51 607.12 1582.27 ;
        RECT  605.52 763.505 607.12 814.27 ;
        RECT  605.52 15.38 607.12 46.27 ;
        RECT  415.52 2299.51 417.12 2352.3 ;
        RECT  415.52 1531.51 417.12 1582.27 ;
        RECT  415.52 763.505 417.12 814.27 ;
        RECT  415.52 15.38 417.12 46.27 ;
        RECT  225.52 2299.53 227.12 2352.3 ;
        RECT  225.52 1531.53 227.12 1579.72 ;
        RECT  225.52 763.53 227.12 811.72 ;
        RECT  225.52 15.38 227.12 43.72 ;
        RECT  35.52 15.38 37.12 2352.3 ;
    END
  END VSS
  OBS
    LAYER Pwell ;
     RECT  0 0 2175 2352.3 ;
    LAYER Nwell ;
     RECT  0 0 2175 2352.3 ;
    LAYER Metal1 ;
     RECT  0 0 2175 2352.3 ;
    LAYER Metal2 ;
     RECT  0 0 2175 2352.3 ;
    LAYER Metal3 ;
     RECT  0 0 2175 2352.3 ;
    LAYER Metal4 ;
     RECT  0 0 2175 2352.3 ;
    LAYER Metal5 ;
        RECT 10 0 2165 34.5 ;
        RECT 10 49.5 2165 79.5 ;
        RECT 10 94.5 2165 124.5 ;
        RECT 10 139.5 2165 169.5 ;
        RECT 10 184.5 2165 214.5 ;
        RECT 10 229.5 2165 259.5 ;
        RECT 10 274.5 2165 304.5 ;
        RECT 10 319.5 2165 349.5 ;
        RECT 10 364.5 2165 394.5 ;
        RECT 10 409.5 2165 439.5 ;
        RECT 10 454.5 2165 484.5 ;
        RECT 10 499.5 2165 529.5 ;
        RECT 10 544.5 2165 574.5 ;
        RECT 10 589.5 2165 619.5 ;
        RECT 10 634.5 2165 664.5 ;
        RECT 10 679.5 2165 709.5 ;
        RECT 10 724.5 2165 754.5 ;
        RECT 10 769.5 2165 799.5 ;
        RECT 10 814.5 2165 844.5 ;
        RECT 10 859.5 2165 889.5 ;
        RECT 10 904.5 2165 934.5 ;
        RECT 10 949.5 2165 979.5 ;
        RECT 10 994.5 2165 1024.5 ;
        RECT 10 1039.5 2165 1069.5 ;
        RECT 10 1084.5 2165 1114.5 ;
        RECT 10 1129.5 2165 1159.5 ;
        RECT 10 1174.5 2165 1204.5 ;
        RECT 10 1219.5 2165 1249.5 ;
        RECT 10 1264.5 2165 1294.5 ;
        RECT 10 1309.5 2165 1339.5 ;
        RECT 10 1354.5 2165 1384.5 ;
        RECT 10 1399.5 2165 1429.5 ;
        RECT 10 1444.5 2165 1474.5 ;
        RECT 10 1489.5 2165 1519.5 ;
        RECT 10 1534.5 2165 1564.5 ;
        RECT 10 1579.5 2165 1609.5 ;
        RECT 10 1624.5 2165 1654.5 ;
        RECT 10 1669.5 2165 1699.5 ;
        RECT 10 1714.5 2165 1744.5 ;
        RECT 10 1759.5 2165 1789.5 ;
        RECT 10 1804.5 2165 1834.5 ;
        RECT 10 1849.5 2165 1879.5 ;
        RECT 10 1894.5 2165 1924.5 ;
        RECT 10 1939.5 2165 1969.5 ;
        RECT 10 1984.5 2165 2014.5 ;
        RECT 10 2029.5 2165 2059.5 ;
        RECT 10 2074.5 2165 2104.5 ;
        RECT 10 2119.5 2165 2149.5 ;
        RECT 10 2164.5 2165 2194.5 ;
        RECT 10 2209.5 2165 2239.5 ;
        RECT 10 2254.5 2165 2284.5 ;
        RECT 10 2299.5 2165 2329.5 ;
  END
END efuse_ctrl
END LIBRARY
